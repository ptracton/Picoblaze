//                              -*- Mode: Verilog -*-
// Filename        : cpu.v
// Description     : Complete Picoblaze Design
// Author          : Philip Tracton
// Created On      : Thu May 21 22:33:37 2015
// Last Modified By: Philip Tracton
// Last Modified On: Thu May 21 22:33:37 2015
// Update Count    : 0
// Status          : Unknown, Use with caution!


module cpu (/*AUTOARG*/ ) ;
 
   
   /*AUTOWIRE*/
   /*AUTOREG*/
endmodule // cpu
